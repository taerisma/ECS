--Auswahlcode für MEP
---------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
---------------------------------
entity MEP is 
	port();
end MEP;
Architecture A1 of MEP is
--Signale
--Konstanten
--Array
begin
end A1;