--SubX
---------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SubX is
	port(
		alpha 	: in std_logic;
		beta	: out std_logic);
end SubX;

architecture Behavioral of SubX is
begin
end Behavioral;