--RAM WbR.vhd