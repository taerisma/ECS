--Auswahlcode für Wein
---------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
---------------------------------
entity Wein is 
	port();
end Wein;
Architecture A1 of Wein is
--Signale
--Konstanten
--Array
begin
end A1;