--SubSubY
-------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SubSubY is
    Port ( 
		x : in  STD_LOGIC;
		y : out  STD_LOGIC);
end SubSubY;

architecture Behavioral of SubSubY is
begin
end Behavioral;