--Auswahlcode für Ferien
---------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
---------------------------------
entity Ferien is 
	port();
end Ferien;
Architecture A1 of Ferien is
--Signale
--Konstanten
--Array
begin
end A1;